`timescale 1ns/1ps
module rv32i_pipeline_regs(); // placeholder file - actual regs in core for clarity
endmodule
